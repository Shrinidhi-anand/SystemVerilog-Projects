// $write("**************************");
// $write("***************************************************\n");  

// $write("**************************");
// $write("***************************************************\n");



//************************GENERATOR**********************//
////filename generator.sv


