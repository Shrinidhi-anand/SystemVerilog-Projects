parameter reg [15:0] ADDR_WIDTH=4;
parameter reg [15:0] DATA_WIDTH=32;
parameter reg [15:0] MEM_SIZE=16;
