
////filename ram_parameter.sv
parameter DATA_WIDTH = 7;
parameter ADDR_WIDTH = 4;
parameter MEM_SIZE = 31;



